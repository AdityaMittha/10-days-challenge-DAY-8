module tb5();reg clk,rst,sin;wire[3:0] pout;sipo uut(clk,rst,sin,pout);initial begin clk=0; forever #5 clk=~clk; end initial begin rst=1; sin=1; #5; rst=0; sin=0; #10; rst=1; sin=1; #10; sin=1; #10; sin=1; #10; sin=0; #10; sin=1; #5; $finish; end endmodule