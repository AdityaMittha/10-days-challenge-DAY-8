module tb9();reg clk,d;wire q;d_flipflop uut(d,clk,q);initial begin clk=0;forever #5 clk=~clk;end initial begin d=0;#10;d=1;#10;d=0;#10;d=1;#10;d=1;#10;d=0;#10;$finish;end endmodule